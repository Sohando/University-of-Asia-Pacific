module _gate(F, A, B);
	input A, B;
	output F;
	and(F, A, B);
endmodule